//--------------------------------------------------------------------------------------------------------------------
// File         : Buffer.sv --> Design of buffer module
// Author       : Manjush Padmamma Venkatesha
// Date Created : March 12 2018
// Description  : Design of Buffer Module, used counter logic to move onto location to location 
//		  either for read or write operation. Data Coherence is handled within the module
//		  Depth is of page size.
//		  Write cant happen from both sides of buffer, either host can write or controller
//		  If one is writing the other could read the same and vice versa.
//		  Once writing of data starts it should write upto complete buffer depth else junk data would be stored on the buffer
//		  Similarly the same happens with read operation
//		  Status signals are asserted once the read operation is completed on both host and controller side
//--------------------------------------------------------------------------------------------------------------------
module Buffer(IBuffer.BufferPorts bufBus);

import BufferDefs :: *;

always_ff @(posedge bufBus.clk) begin				//for buffer to host interface opeartion
	if(bufBus.buf_sel && host_addr < Buf_Depth) begin
		bufBus.host_buf_status <= 0;
		if(bufBus.buf_we && !bufBus.buf_cntrl_status && !buf_write_flag) begin  //buffer write opeartion on host side
			buf_mem[host_addr] <= bufBus.buf_in;
			host_addr <= host_addr + 1;
			cntrl_read_flag <= 1;
		end	
		else
			host_addr <= 0;

		if(bufBus.buf_re && buf_read_flag) begin	//buffer read opeartion on host side
			bufBus.buf_out <= buf_mem[host_addr];
			host_addr <= host_addr + 1;
		end
		if(host_addr == Buf_Depth - 1) begin		//controlling status on host read operation
			if(buf_read_flag)
				bufBus.host_buf_status <= 1;
			else
				bufBus.host_buf_status <= 0;
		end
	end
	else if(host_addr == Buf_Depth) begin			//when buffer depth is reached 
		if(bufBus.buf_sel) begin			//avoid overwrite and over
			if(bufBus.buf_re) begin
				$display("read from buffer to host completed!!!! dont read for more @%0d",$time);
			end
			if(bufBus.buf_we) begin
				buf_write_flag <=1;
				$display("write from host to buffer--> buffer full @%0d",$time);
			end
		end
		
		bufBus.host_buf_status <= 0;
		cntrl_write_flag <= 0;				//reset all flags once it is hovered througout buffer depth
		buf_read_flag <= 0;
		host_addr <= 0;
	end
	else begin						//reset address and status once buffer is idle or operation is completed
		host_addr <= 0;
		bufBus.host_buf_status <= 0;
	end

	if(bufBus.cntrl_sel && cntrl_addr < Buf_Depth) begin	//for buffer to controller interface operation
		bufBus.buf_cntrl_status <= 0;
		if(bufBus.cntrl_re && cntrl_read_flag) begin	//buffer read operation on controller side
			bufBus.cntrl_out <= buf_mem[cntrl_addr];
			cntrl_addr <= cntrl_addr + 1;
		end

		if(bufBus.cntrl_we && !bufBus.host_buf_status && !cntrl_write_flag) begin	//buffer write operation on controller side
			buf_mem[cntrl_addr] <= bufBus.cntrl_in;

			cntrl_addr <= cntrl_addr + 1;
			buf_read_flag <= 1;
		end
		if(cntrl_addr == Buf_Depth - 1) begin		//controlling status on controller read operation
			if(cntrl_read_flag)
				bufBus.buf_cntrl_status <= 1;
			else
				bufBus.buf_cntrl_status <= 0;
		end
	end
	else if(cntrl_addr == Buf_Depth) begin			//when buffer depth is reached 
		if (bufBus.cntrl_sel) begin			//avoid overwrite and over read of data
			if(bufBus.cntrl_re) begin
				$display("read from buffer to controller completed!!!! dont read for more @%0d",$time);
			end
			if(bufBus.cntrl_we) begin
				cntrl_write_flag <= 1;
				$display("write from controller to buffer--> buffer full @%0d",$time);
			end
		end
		bufBus.buf_cntrl_status <= 0;
		buf_write_flag <= 0;				//reset all flags once it is hovered
		cntrl_read_flag <= 0;
		cntrl_addr <= 0;
	end
	else begin						//reset address and status once buffer is idle or operation is completed
		cntrl_addr <= 0;
		bufBus.buf_cntrl_status <= 0;
	end
	
end
endmodule : Buffer
